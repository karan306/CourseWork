--
-- Copyright (C) 2009-2012 Chris McClelland
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU Lesser General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity top_level is
	port(
		-- FX2LP interface ---------------------------------------------------------------------------
		sys_clk			: in 	  std_logic;
		fx2Clk_in      : in    std_logic;                    -- 48MHz clock from FX2LP
		fx2Addr_out    : out   std_logic_vector(1 downto 0); -- select FIFO: "00" for EP2OUT, "10" for EP6IN
		fx2Data_io     : inout std_logic_vector(7 downto 0); -- 8-bit data to/from FX2LP

		-- When EP2OUT selected:
		fx2Read_out    : out   std_logic;                    -- asserted (active-low) when reading from FX2LP
		fx2OE_out      : out   std_logic;                    -- asserted (active-low) to tell FX2LP to drive bus
		fx2GotData_in  : in    std_logic;                    -- asserted (active-high) when FX2LP has data for us

		-- When EP6IN selected:
		fx2Write_out   : out   std_logic;                    -- asserted (active-low) when writing to FX2LP
		fx2GotRoom_in  : in    std_logic;                    -- asserted (active-high) when FX2LP has room for more data from us
		fx2PktEnd_out  : out   std_logic;                    -- asserted (active-low) when a host read needs to be committed early

		-- Onboard peripherals -----------------------------------------------------------------------
		--sseg_out       : out   std_logic_vector(7 downto 0); -- seven-segment display cathodes (one for each segment)
		--anode_out      : out   std_logic_vector(3 downto 0); -- seven-segment display anodes (one for each digit)
		led_out        : out   std_logic_vector(7 downto 0); -- eight LEDs
		sw_in          : in    std_logic_vector(7 downto 0);  -- eight switches
		reset 	      : in	  std_logic;
		left	 	      : in	  std_logic;
		right 	      : in	  std_logic;
		up		 	      : in	  std_logic;
		down	 	      : in	  std_logic;
		-------------------------------------------------------------------------------------------------------------------------
		uart_rx	: in std_logic;
		uart_tx	: out std_logic
	);
end entity;

architecture structural of top_level is
	-- Channel read/write interface -----------------------------------------------------------------
	signal chanAddr  : std_logic_vector(6 downto 0);  -- the selected channel (0-127)

	-- Host >> FPGA pipe:
	signal h2fData   : std_logic_vector(7 downto 0);  -- data lines used when the host writes to a channel
	signal h2fValid  : std_logic;                     -- '1' means "on the next clock rising edge, please accept the data on h2fData"
	signal h2fReady  : std_logic;                     -- channel logic can drive this low to say "I'm not ready for more data yet"

	-- Host << FPGA pipe:
	signal f2hData   : std_logic_vector(7 downto 0);  -- data lines used when the host reads from a channel
	signal f2hValid  : std_logic;                     -- channel logic can drive this low to say "I don't have data ready for you"
	signal f2hReady  : std_logic;     					  -- '1' means "on the next clock rising edge, put your next byte of data on f2hData"
	-- ----------------------------------------------------------------------------------------------
	

	-- Needed so that the comm_fpga_fx2 module can drive both fx2Read_out and fx2OE_out
	signal fx2Read   : std_logic;

	-- Reset signal so host can delay startup
	signal fx2Reset  : std_logic;
	
	--------------------------------------------------------------------------------------------------------
	
	signal left_b	  : std_logic;
	signal right_b	  : std_logic;
	signal up_b	 	  : std_logic;
	signal down_b	  : std_logic;
	
	signal	wr_en  :  std_logic; --20102016
	signal 	rd_en  :  std_logic; --20102016
	signal	full   :  std_logic; --20102016
	signal	empty  :  std_logic; --20102016);
	signal 	start	 :  std_logic;
	signal 	pop	 :  std_logic;
	signal 	data_out	 :  std_logic_vector(7 downto 0);
	
	component debouncer
        port(clk: in STD_LOGIC;
            button: in STD_LOGIC;
            button_deb: out STD_LOGIC);
   end component;
	 
	 component uart is
		port (clk 	 : in std_logic;
				rst 	 : in std_logic;
				rx	 	 : in std_logic;
				tx	 	 : out std_logic;
				data_in	 : in std_logic_vector(7 downto 0);
				data_out	 : out std_logic_vector(7 downto 0);
				pop 	 : in std_logic;
				start	 : in std_logic;
				--Signals pulled on Atlys LEDs for debugging
				Bwr_en  : out std_logic; --20102016
				Brd_en  : out std_logic; --20102016
				Bfull   : out std_logic;--20102016
				Bempty  : out std_logic); --20102016
	 end component uart;	


begin
		
	i_uart : uart port map (pop=>pop,data_in=>sw_in,data_out=>data_out,start=>start,clk => sys_clk, rst => reset, rx => uart_rx, tx => uart_tx, Bwr_en => wr_en, Brd_en => rd_en, Bfull => full, Bempty => empty);  --20102016
	
	-- CommFPGA module
	fx2Read_out <= fx2Read;
	fx2OE_out <= fx2Read;
	fx2Addr_out(0) <=  -- So fx2Addr_out(1)='0' selects EP2OUT, fx2Addr_out(1)='1' selects EP6IN
		'0' when fx2Reset = '0'
		else 'Z';
	comm_fpga_fx2 : entity work.comm_fpga_fx2
		port map(
			clk_in         => fx2Clk_in,
			reset_in       => '0',
			reset_out      => fx2Reset,
			
			-- FX2LP interface
			fx2FifoSel_out => fx2Addr_out(1),
			fx2Data_io     => fx2Data_io,
			fx2Read_out    => fx2Read,
			fx2GotData_in  => fx2GotData_in,
			fx2Write_out   => fx2Write_out,
			fx2GotRoom_in  => fx2GotRoom_in,
			fx2PktEnd_out  => fx2PktEnd_out,

			-- DVR interface -> Connects to application module
			chanAddr_out   => chanAddr,
			h2fData_out    => h2fData,
			h2fValid_out   => h2fValid,
			h2fReady_in    => h2fReady,
			f2hData_in     => f2hData,
			f2hValid_in    => f2hValid,
			f2hReady_out   => f2hReady
		);
		
		debouncer1: debouncer
              port map (clk => fx2Clk_in,
                        button => left,
                        button_deb => left_b);

		debouncer2: debouncer
						  port map (clk => fx2Clk_in,
										button => right,
										button_deb => right_b);

		debouncer3: debouncer
						  port map (clk => fx2Clk_in,
										button => up,
										button_deb => up_b);

		debouncer4: debouncer
						  port map (clk => fx2Clk_in,
										button => down,
										button_deb => down_b);

	-- Switches & LEDs application
	swled_app : entity work.swled
		port map(
			clk_in       => fx2Clk_in,
			reset_in     => reset,
			-- DVR interface -> Connects to comm_fpga module
			chanAddr_in  => chanAddr,
			h2fData_in   => h2fData,
			h2fValid_in  => h2fValid,
			h2fReady_out => h2fReady,
			f2hData_out  => f2hData,
			f2hValid_out => f2hValid,
			f2hReady_in  => f2hReady,
			
			-- External interface
			--sseg_out     => sseg_out,
			--anode_out    => anode_out,
			led_out      => led_out,
			sw_in        => sw_in,
			left				=> left_b,
			right				=> right_b,
			up					=> up_b,
			down				=> down_b,
			empty				=> empty,
			start				=>start,
			data				=>data_out,
			pop				=>pop
		);
end architecture;
